library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.INTEGER_VECTOR.all;


ENTITY VGA IS
GENERIC (
	ALIEN_NUMBER : INTEGER RANGE -10 TO 1200 := 32;
	SHOTS_NUMBER : INTEGER RANGE -10 TO 1200 := 10;
	SHOT_SIZE_X : INTEGER RANGE -10 TO 1200 := 10;
	SHOT_SIZE_Y : INTEGER RANGE -10 TO 1200 := 40;
	BATTLEFIELD_SIZE : INTEGER RANGE -10 TO 1200 := 900;
	INITIAL_PLAYER_LIVES : INTEGER RANGE -10 TO 1200 := 3;
	NUMBER_OF_LEVELS : INTEGER RANGE -10 TO 1200 := 3
);
PORT(
	CLOCK_50: IN STD_LOGIc;
	GAME_STATUS: IN INTEGER RANGE 0 TO 3;
	LEVEL : IN INTEGER RANGE 0 TO NUMBER_OF_LEVELS;
	LIVES_P1: IN INTEGER RANGE 0 TO INITIAL_PLAYER_LIVES;
	LIVES_P2: IN INTEGER RANGE 0 TO INITIAL_PLAYER_LIVES;
	SCORE: IN INTEGER RANGE -10 TO 1200;
	ENEMY_SHIPS_X : IN INTEGER_VECTOR(ALIEN_NUMBER-1 downto 0);
	ENEMY_SHIPS_Y : IN INTEGER_VECTOR(ALIEN_NUMBER-1 downto 0);
	ENEMY_SHOTS_X : IN INTEGER_VECTOR(SHOTS_NUMBER-1 downto 0);
	ENEMY_SHOTS_Y : IN INTEGER_VECTOR(SHOTS_NUMBER-1 downto 0);
	SHOT_X_P1 : IN INTEGER RANGE -10 TO 1200;
	SHOT_Y_P1 : IN INTEGER RANGE -10 TO 1200;
	SHOT_X_P2 : IN INTEGER RANGE -10 TO 1200;
	SHOT_Y_P2 : IN INTEGER RANGE -10 TO 1200;
	SHIP_X_P1 : IN INTEGER RANGE -10 TO 1200;
	SHIP_Y_P1 : IN INTEGER RANGE -10 TO 1200;
	SHIP_X_P2 : IN INTEGER RANGE -10 TO 1200;
	SHIP_Y_P2 : IN INTEGER RANGE -10 TO 1200;
	VGA_HS,VGA_VS:OUT STD_LOGIC;
	VGA_R,VGA_B,VGA_G: OUT STD_LOGIC_VECTOR(3 downto 0)
);
END VGA;


ARCHITECTURE MAIN OF VGA IS
SIGNAL VGACLK:STD_LOGIC;
SIGNAL RESET:STD_LOGIC := '0';

	COMPONENT SYNC IS
		GENERIC (
			ALIEN_NUMBER : INTEGER RANGE -10 TO 1200 := 32;
			SHOTS_NUMBER : INTEGER RANGE -10 TO 1200 := 10;
			SHOT_SIZE_X : INTEGER RANGE -10 TO 1200 := 10;
			SHOT_SIZE_Y : INTEGER RANGE -10 TO 1200 := 40;
			BATTLEFIELD_SIZE : INTEGER RANGE -10 TO 1200 := 900
		);
		PORT(
			CLK: IN STD_LOGIC;
			HSYNC: OUT STD_LOGIC;
			VSYNC: OUT STD_LOGIC;
			GAME_STATUS: IN INTEGER RANGE 0 TO 3;
			LEVEL : IN INTEGER RANGE 0 TO 7;
			LIVES_P1: IN INTEGER RANGE 0 TO 3;
			LIVES_P2: IN INTEGER RANGE 0 TO 3;
			SCORE: IN INTEGER RANGE -10 TO 1200;
			ENEMY_SHIPS_X : IN INTEGER_VECTOR(ALIEN_NUMBER-1 downto 0);
			ENEMY_SHIPS_Y : IN INTEGER_VECTOR(ALIEN_NUMBER-1 downto 0);
			ENEMY_SHOTS_X : IN INTEGER_VECTOR(SHOTS_NUMBER-1 downto 0);
			ENEMY_SHOTS_Y : IN INTEGER_VECTOR(SHOTS_NUMBER-1 downto 0);
			SHOT_X_P1 : IN INTEGER RANGE 0 TO 1200;
			SHOT_Y_P1 : IN INTEGER RANGE 0 TO 1200;
			SHOT_X_P2 : IN INTEGER RANGE 0 TO 1200;
			SHOT_Y_P2 : IN INTEGER RANGE 0 TO 1200;
			SHIP_X_P1 : IN INTEGER RANGE 0 TO 1200;
			SHIP_Y_P1 : IN INTEGER RANGE 0 TO 1200;
			SHIP_X_P2 : IN INTEGER RANGE 0 TO 1200;
			SHIP_Y_P2 : IN INTEGER RANGE 0 TO 1200;
			R: OUT STD_LOGIC_VECTOR(3 downto 0);
			G: OUT STD_LOGIC_VECTOR(3 downto 0);
			B: OUT STD_LOGIC_VECTOR(3 downto 0)
		);
	END COMPONENT SYNC;

	component pll is
		port (
			clk_out_clk : out std_logic;        -- clk
			clk_in_clk  : in  std_logic := 'X'; -- clk
			reset_reset  : in  std_logic := 'X'  -- reset
		);
	END COMPONENT pll;
	 
 BEGIN
 
 C: pll PORT MAP (VGACLK,CLOCK_50,RESET);
 C1: SYNC generic map (
					ALIEN_NUMBER => ALIEN_NUMBER,
					SHOTS_NUMBER => SHOTS_NUMBER,
					SHOT_SIZE_X => SHOT_SIZE_X,
					SHOT_SIZE_Y => SHOT_SIZE_Y,
					BATTLEFIELD_SIZE => BATTLEFIELD_SIZE
				) 
				PORT MAP(VGACLK,VGA_HS,VGA_VS,GAME_STATUS,LEVEL,LIVES_P1,LIVES_P2,SCORE,
						 ENEMY_SHIPS_X,ENEMY_SHIPS_Y,ENEMY_SHOTS_X,ENEMY_SHOTS_Y,SHOT_X_P1,SHOT_Y_P1,
						 SHOT_X_P2,SHOT_Y_P2,SHIP_X_P1,SHIP_Y_P1, SHIP_X_P2,SHIP_Y_P2,VGA_R,VGA_G,VGA_B);
 
 END MAIN;
 